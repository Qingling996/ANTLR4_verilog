/* 区块注释【可能有可能没有】 */
// 单行注释【可能有可能没有】

// 与编译指令【可能有可能没有】
`timescale 1ns/1ns
`define hello 25
// `include "VerilogLexer.g4"

module module_name 
    #(
        // 可能存在的端口参数
    )
    (
        // 端口声明
        // input [wire] [signed] [range] 端口名，
        // output [wire | reg] [signed] [range] 端口名，
        // inout [wire] [signed] [range] 端口名，
    );

/* ================================================================================================  */
/*                                              信号声明                                              */
/* ================================================================================================  */
// (parameter | localparam) [signed] [range] 参数名;
// reg  [signed] [range] 变量名;
reg      [03:00]        S_add; //
// wire [signed] [range] 变量名;
// integer 变量名;
// real 变量名;
// time 变量名;

/* ================================================================================================  */
/*                                             模块实例化                                             */
/* ================================================================================================  */

/* ================================================================================================  */
/*                                          连续赋值和过程块                                          */
/* ================================================================================================  */
// assign 信号名 = 表达式;

// always /* @(敏感信号列表) */  
    // statement

// initial
    // statement
initial begin 
    case(S_add)
        2:S_add <= 3;
        default: ;
    endcase
    if(S_add)begin
        
    end
end 
/* ================================================================================================  */
/*                                          任务/函数/生成块                                          */
/* ================================================================================================  */
// task
    // statement

// function
    // statement

// generate
    // statement

/* ================================================================================================  */
/*                                                                                                  */
/* ================================================================================================  */

/* statement
    1、循环
    2、条件 (if - else if - else)
    3、条件 (case/casez/casex)
    4、
    ｝ 
*/

endmodule 


